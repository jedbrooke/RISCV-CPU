`timescale 1ns / 100ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/14/2020 12:17:55 PM
// Design Name: 
// Module Name: add_and_subtract_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module add_and_subtract_tb(

    );
    parameter WIDTH = 32;

    reg [WIDTH-1:0] a;
    reg [WIDTH-1:0] b;
    wire cout;
    wire [WIDTH-1:0] sum;
    reg subtract;
    wire add_correct;
    wire sub_correct;
    
    add_and_subtract uut(.a(a), .b(b), .cout(cout), .sum(sum), .subtract(subtract) );
    
    assign add_correct = (subtract ? (a - b) : (a + b)) == sum;

    
    initial begin
        a = 1;
        b = 1;
        subtract = 0;
        a = 3175089953;
        b = 3973635537;
        #5;
        a = 655546290;
        b = 2720499003;
        #5;
        a = 710837918;
        b = 1558857175;
        #5;
        a = 201962729;
        b = 4289023901;
        #5;
        a = 642745811;
        b = 3580119396;
        #5;
        a = 2576462504;
        b = 4144025494;
        #5;
        a = 4054230487;
        b = 1113334425;
        #5;
        a = 46302133;
        b = 2948875240;
        #5;
        a = 2400551831;
        b = 2045140421;
        #5;
        a = 1625835701;
        b = 4130241201;
        #5;
        a = 2220213121;
        b = 4212933799;
        #5;
        a = 1729996874;
        b = 680139810;
        #5;
        a = 550986017;
        b = 2059669277;
        #5;
        a = 2800386767;
        b = 2705563037;
        #5;
        a = 3495277561;
        b = 1023943478;
        #5;
        a = 3443447381;
        b = 770601583;
        #5;
        a = 3286513444;
        b = 1761934228;
        #5;
        a = 452077134;
        b = 1592047779;
        #5;
        a = 3932792380;
        b = 3805019076;
        #5;
        a = 2701214133;
        b = 1556581075;
        #5;
        a = 992050908;
        b = 3765308988;
        #5;
        a = 1420327208;
        b = 2450508766;
        #5;
        a = 3824615452;
        b = 3680597417;
        #5;
        a = 2909093241;
        b = 2632534260;
        #5;
        a = 3139530764;
        b = 2738760048;
        #5;
        a = 1505590233;
        b = 3806682887;
        #5;
        a = 1834032090;
        b = 2189943533;
        #5;
        a = 1824487651;
        b = 125197716;
        #5;
        a = 3900123347;
        b = 540356755;
        #5;
        a = 3504427652;
        b = 1830360565;
        #5;
        a = 3420017261;
        b = 3593165175;
        #5;
        a = 3518633926;
        b = 4109194362;
        #5;
        a = 3713101738;
        b = 1465849377;
        #5;
        a = 3270366286;
        b = 1396227371;
        #5;
        a = 3193070586;
        b = 3980903974;
        #5;
        a = 3687939697;
        b = 2642171907;
        #5;
        a = 919560273;
        b = 2279923163;
        #5;
        a = 2161889683;
        b = 1277490992;
        #5;
        a = 1619412412;
        b = 1938412132;
        #5;
        a = 144220104;
        b = 3239581909;
        #5;
        a = 2808251350;
        b = 4101588556;
        #5;
        a = 604406880;
        b = 2905376522;
        #5;
        a = 1429047094;
        b = 1240986476;
        #5;
        a = 1885367279;
        b = 1641511314;
        #5;
        a = 512150999;
        b = 3229760740;
        #5;
        a = 3712450854;
        b = 3866697716;
        #5;
        a = 480842645;
        b = 3699097690;
        #5;
        a = 1742516274;
        b = 3227518876;
        #5;
        a = 3725438249;
        b = 3882464847;
        #5;
        a = 2138723706;
        b = 4071033972;
        #5;
        a = 798203518;
        b = 881487960;
        #5;
        a = 248188881;
        b = 66652665;
        #5;
        a = 3494115148;
        b = 3347461814;
        #5;
        a = 3284593429;
        b = 2087022174;
        #5;
        a = 2632560601;
        b = 2307773265;
        #5;
        a = 2659708416;
        b = 354430149;
        #5;
        a = 515715565;
        b = 4038917392;
        #5;
        a = 3259723620;
        b = 1027244646;
        #5;
        a = 2863940321;
        b = 285485002;
        #5;
        a = 3960595462;
        b = 2344345715;
        #5;
        a = 2906877957;
        b = 2844045726;
        #5;
        a = 3858206388;
        b = 2663504094;
        #5;
        a = 1527929944;
        b = 873974887;
        #5;
        a = 1577082492;
        b = 3296861250;
        #5;
        a = 3750759199;
        b = 3950070922;
        #5;
        a = 3601096783;
        b = 2443022716;
        #5;
        a = 3837017414;
        b = 1985592349;
        #5;
        a = 1520171210;
        b = 3745958848;
        #5;
        a = 3668585424;
        b = 908971079;
        #5;
        a = 1891151759;
        b = 3937700836;
        #5;
        a = 2777373840;
        b = 2977612351;
        #5;
        a = 741750576;
        b = 1259871975;
        #5;
        a = 344400613;
        b = 4069396920;
        #5;
        a = 3875176686;
        b = 3313813968;
        #5;
        a = 1065623479;
        b = 2999093055;
        #5;
        a = 533888253;
        b = 2772846242;
        #5;
        a = 299516215;
        b = 855652016;
        #5;
        a = 27106328;
        b = 1653938094;
        #5;
        a = 2908129109;
        b = 1915601595;
        #5;
        a = 1067761780;
        b = 45973596;
        #5;
        a = 2820614285;
        b = 516867084;
        #5;
        a = 1793472547;
        b = 2377659629;
        #5;
        a = 3603228096;
        b = 1529753954;
        #5;
        a = 659149349;
        b = 2607415163;
        #5;
        a = 3885954908;
        b = 3024335716;
        #5;
        a = 928509347;
        b = 2954304352;
        #5;
        a = 3755245380;
        b = 4285425757;
        #5;
        a = 3176980379;
        b = 2145439323;
        #5;
        a = 2651106366;
        b = 3783939605;
        #5;
        a = 3907676297;
        b = 3305326779;
        #5;
        a = 2891764430;
        b = 4039022565;
        #5;
        a = 1623297122;
        b = 2256336357;
        #5;
        a = 3594944361;
        b = 2540585454;
        #5;
        a = 2223372635;
        b = 1953139727;
        #5;
        a = 705473006;
        b = 3358280543;
        #5;
        a = 2781547581;
        b = 1471694508;
        #5;
        a = 3418634363;
        b = 3325262049;
        #5;
        a = 684380777;
        b = 3687399393;
        #5;
        a = 2726558086;
        b = 2435191187;
        #5;
        a = 3340168906;
        b = 4084575728;
        #5;
        $finish;
    end
//    always begin
//        #5 a = a << 1;
//    end
    
//    always @(negedge a[WIDTH-1]) begin
//        b = b << 1;
//        a = 1;
//    end
    
//    always @* begin
//        if(b[WIDTH - 1]) begin
//            $finish;
//        end
//    end
    
    
    
endmodule
